module main

fn main() {
	eprintln('Update disabled.')
	exit(1)
}
